//==================================================
// Author : Chris Le
// Email  : lehoangcuong1990@gmail.com
// Date   : July 08, 2018
//==================================================
 
`ifndef _ALU_REG_PREDICTOR_
`define _ALU_REG_PREDICTOR_
typedef uvm_reg_predictor#(apb_seq_item) alu_reg_predictor;
`endif
