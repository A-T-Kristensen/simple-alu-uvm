//==================================================
// Author : Chris Le
// Email  : lehoangcuong1990@gmail.com
// Date   : July 08, 2018
//==================================================
 
`ifndef _ALU_SEQR_
`define _ALU_SEQR_
typedef uvm_sequencer#(alu_trans) alu_seqr;
`endif
